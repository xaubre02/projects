-- IVH project, Vojtech Mrazek, xmraze06
-- Vraci dekodovani znaku 8x16 podle vstupu
-- 
library IEEE;
use IEEE.std_logic_1164.ALL;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity char_rom is
	Generic (
		SIZE : integer := 4
	);
	Port (
		ADDRESS : in std_logic_vector(SIZE-1 downto 0);
		ROW : in std_logic_vector(3 downto 0);
		COLUMN : in std_logic_vector(2 downto 0);
		DATA : out std_logic
	);
end char_rom;

architecture behv of char_rom is
	type t_mem is array (0 to (2**SIZE)-1) of std_logic_vector(0 to 127);
	constant rommem : t_mem :=(
--znak  => "   1   |   2   |   3   |   4   |   5   |   6   |   7   |   8   |   9   |  10   |   11  |   12  |  13   |   14  |   15  |   16  |)
		 0 => "00000000000000000000000000000000000000000001110000100010001000100010001000100010001000100001110000000000000000000000000000000000", -- 0
		 1 => "00000000000000000000000000000000000000000011111000001000000010000000100000001000000010000000110000000000000000000000000000000000", -- 1
		 2 => "00000000000000000000000000000000000000000011111000000010000001000000100000010000001000100001110000000000000000000000000000000000", -- 2
		 3 => "00000000000000000000000000000000000000000001110000100010001000000001100000100000001000100001110000000000000000000000000000000000", -- 3
		 4 => "00000000000000000000000000000000000000000011100000010000001111100001001000010100000110000001000000000000000000000000000000000000", -- 4
		 5 => "00000000000000000000000000000000000000000001110000100010001000000001110000000100000001000011110000000000000000000000000000000000", -- 5
		 6 => "00000000000000000000000000000000000000000001110000100010001000100001111000000010000001000011100000000000000000000000000000000000", -- 6
		 7 => "00000000000000000000000000000000000000000000100000001000000100000001000000100000001000100011111000000000000000000000000000000000", -- 7
		 8 => "00000000000000000000000000000000000000000001110000100010001000100001110000100010001000100001110000000000000000000000000000000000", -- 8
		 9 => "00000000000000000000000000000000000000000000111000010000001000000011110000100010001000100001110000000000000000000000000000000000", -- 9
		--10 => "00000000000000000000000000000000000000000111011100100010000111000001010000010100000010000000110000000000000000000000000000000000", -- A
	 	--11 => "00000000000000000000000000000000000000000001111100100010001000100001111000100010001000100001111100000000000000000000000000000000", -- B
		--12 => "00000000000000000000000000000000000000000001110000100010000000100000001000000010001000100011110000000000000000000000000000000000", -- C
		--13 => "00000000000000000000000000000000000000000000111100010010001000100010001000100010000100100000111100000000000000000000000000000000", -- D
		--14 => "00000000000000000000000000000000000000000011111000100100000101000001110000010100001001000011111000000000000000000000000000000000", -- E
		--15 => "00000000000000000000000000000000000000000000111000000100000101000001110000010100001001000011111000000000000000000000000000000000", -- F
					 
		 others => (others=>'-') -- others don't care
		); 
	
begin
	vyhodnoceni: process (ADDRESS, ROW, COLUMN) is 
   	variable var_data : std_logic_vector(127 downto 0);
	begin
		var_data := rommem(conv_integer(ADDRESS));
		data <= var_data(conv_integer(ROW & COLUMN));
      
	end process vyhodnoceni;
 
end behv;
